e(1,2).
e(2,3).
e(1,3).
path(X,Y):-e(X,Y).
path(X,Y):-path(X,Z),path(Z,Y).